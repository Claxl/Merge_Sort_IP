
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "df_fifo_interface.svh"
`include "df_fifo_monitor.svh"
`include "df_process_interface.svh"
`include "df_process_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);

    df_fifo_intf fifo_intf_1(clock,reset);
    assign fifo_intf_1.rd_en = AESL_inst_merge_sort.output_r_c_U.if_read & AESL_inst_merge_sort.output_r_c_U.if_empty_n;
    assign fifo_intf_1.wr_en = AESL_inst_merge_sort.output_r_c_U.if_write & AESL_inst_merge_sort.output_r_c_U.if_full_n;
    assign fifo_intf_1.fifo_rd_block = ~(AESL_inst_merge_sort.write_output_U0.output_r_blk_n);
    assign fifo_intf_1.fifo_wr_block = ~(AESL_inst_merge_sort.entry_proc_U0.output_r_c_blk_n);
    assign fifo_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_1;
    csv_file_dump cstatus_csv_dumper_1;
    df_fifo_monitor fifo_monitor_1;
    df_fifo_intf fifo_intf_2(clock,reset);
    assign fifo_intf_2.rd_en = AESL_inst_merge_sort.left_stream_U.if_read & AESL_inst_merge_sort.left_stream_U.if_empty_n;
    assign fifo_intf_2.wr_en = AESL_inst_merge_sort.left_stream_U.if_write & AESL_inst_merge_sort.left_stream_U.if_full_n;
    assign fifo_intf_2.fifo_rd_block = ~(AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.left_stream_blk_n);
    assign fifo_intf_2.fifo_wr_block = ~(AESL_inst_merge_sort.read_input_U0.left_stream_blk_n);
    assign fifo_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_2;
    csv_file_dump cstatus_csv_dumper_2;
    df_fifo_monitor fifo_monitor_2;
    df_fifo_intf fifo_intf_3(clock,reset);
    assign fifo_intf_3.rd_en = AESL_inst_merge_sort.right_stream_U.if_read & AESL_inst_merge_sort.right_stream_U.if_empty_n;
    assign fifo_intf_3.wr_en = AESL_inst_merge_sort.right_stream_U.if_write & AESL_inst_merge_sort.right_stream_U.if_full_n;
    assign fifo_intf_3.fifo_rd_block = ~(AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.right_stream_blk_n);
    assign fifo_intf_3.fifo_wr_block = ~(AESL_inst_merge_sort.read_input_3_U0.right_stream_blk_n);
    assign fifo_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_3;
    csv_file_dump cstatus_csv_dumper_3;
    df_fifo_monitor fifo_monitor_3;
    df_fifo_intf fifo_intf_4(clock,reset);
    assign fifo_intf_4.rd_en = AESL_inst_merge_sort.tmp_left_U.if_read & AESL_inst_merge_sort.tmp_left_U.if_empty_n;
    assign fifo_intf_4.wr_en = AESL_inst_merge_sort.tmp_left_U.if_write & AESL_inst_merge_sort.tmp_left_U.if_full_n;
    assign fifo_intf_4.fifo_rd_block = ~(AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.tmp_left_blk_n);
    assign fifo_intf_4.fifo_wr_block = ~(AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.tmp_left_blk_n);
    assign fifo_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_4;
    csv_file_dump cstatus_csv_dumper_4;
    df_fifo_monitor fifo_monitor_4;
    df_fifo_intf fifo_intf_5(clock,reset);
    assign fifo_intf_5.rd_en = AESL_inst_merge_sort.tmp_right_U.if_read & AESL_inst_merge_sort.tmp_right_U.if_empty_n;
    assign fifo_intf_5.wr_en = AESL_inst_merge_sort.tmp_right_U.if_write & AESL_inst_merge_sort.tmp_right_U.if_full_n;
    assign fifo_intf_5.fifo_rd_block = ~(AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.tmp_right_blk_n);
    assign fifo_intf_5.fifo_wr_block = ~(AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.tmp_right_blk_n);
    assign fifo_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_5;
    csv_file_dump cstatus_csv_dumper_5;
    df_fifo_monitor fifo_monitor_5;
    df_fifo_intf fifo_intf_6(clock,reset);
    assign fifo_intf_6.rd_en = AESL_inst_merge_sort.tmp_U.if_read & AESL_inst_merge_sort.tmp_U.if_empty_n;
    assign fifo_intf_6.wr_en = AESL_inst_merge_sort.tmp_U.if_write & AESL_inst_merge_sort.tmp_U.if_full_n;
    assign fifo_intf_6.fifo_rd_block = ~(AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.tmp_blk_n);
    assign fifo_intf_6.fifo_wr_block = ~(AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.tmp_blk_n & AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.tmp_blk_n);
    assign fifo_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_6;
    csv_file_dump cstatus_csv_dumper_6;
    df_fifo_monitor fifo_monitor_6;
    df_fifo_intf fifo_intf_7(clock,reset);
    assign fifo_intf_7.rd_en = AESL_inst_merge_sort.output_stream_U.if_read & AESL_inst_merge_sort.output_stream_U.if_empty_n;
    assign fifo_intf_7.wr_en = AESL_inst_merge_sort.output_stream_U.if_write & AESL_inst_merge_sort.output_stream_U.if_full_n;
    assign fifo_intf_7.fifo_rd_block = ~(AESL_inst_merge_sort.write_output_U0.output_stream_blk_n);
    assign fifo_intf_7.fifo_wr_block = ~(AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.output_stream_blk_n);
    assign fifo_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_7;
    csv_file_dump cstatus_csv_dumper_7;
    df_fifo_monitor fifo_monitor_7;

logic region_0_idle;
logic [31:0] region_0_start_cnt;
logic [31:0] region_0_done_cnt;
assign region_0_idle = (region_0_start_cnt == region_0_done_cnt) && AESL_inst_merge_sort.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_start_cnt <= 32'h0;
    else if (AESL_inst_merge_sort.ap_start == 1'b1 && AESL_inst_merge_sort.ap_ready == 1'b1)
        region_0_start_cnt <= region_0_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_done_cnt <= 32'h0;
    else if (AESL_inst_merge_sort.ap_done == 1'b1)
        region_0_done_cnt <= region_0_done_cnt + 32'h1;
    else;
end


    df_process_intf process_intf_1(clock,reset);
    assign process_intf_1.ap_start = AESL_inst_merge_sort.entry_proc_U0.ap_start;
    assign process_intf_1.ap_ready = AESL_inst_merge_sort.entry_proc_U0.ap_ready;
    assign process_intf_1.ap_done = AESL_inst_merge_sort.entry_proc_U0.ap_done;
    assign process_intf_1.ap_continue = AESL_inst_merge_sort.entry_proc_U0.ap_continue;
    assign process_intf_1.real_start = AESL_inst_merge_sort.entry_proc_U0.real_start;
    assign process_intf_1.pin_stall = 1'b0;
    assign process_intf_1.pout_stall = 1'b0 | ~AESL_inst_merge_sort.entry_proc_U0.output_r_c_blk_n;
    assign process_intf_1.cin_stall = 1'b0;
    assign process_intf_1.cout_stall = 1'b0;
    assign process_intf_1.region_idle = region_0_idle;
    assign process_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_1;
    csv_file_dump pstatus_csv_dumper_1;
    df_process_monitor process_monitor_1;
    df_process_intf process_intf_2(clock,reset);
    assign process_intf_2.ap_start = AESL_inst_merge_sort.read_input_U0.ap_start;
    assign process_intf_2.ap_ready = AESL_inst_merge_sort.read_input_U0.ap_ready;
    assign process_intf_2.ap_done = AESL_inst_merge_sort.read_input_U0.ap_done;
    assign process_intf_2.ap_continue = AESL_inst_merge_sort.read_input_U0.ap_continue;
    assign process_intf_2.real_start = AESL_inst_merge_sort.read_input_U0.real_start;
    assign process_intf_2.pin_stall = 1'b0;
    assign process_intf_2.pout_stall = 1'b0 | ~AESL_inst_merge_sort.read_input_U0.left_stream_blk_n;
    assign process_intf_2.cin_stall = 1'b0;
    assign process_intf_2.cout_stall = 1'b0;
    assign process_intf_2.region_idle = region_0_idle;
    assign process_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_2;
    csv_file_dump pstatus_csv_dumper_2;
    df_process_monitor process_monitor_2;
    df_process_intf process_intf_3(clock,reset);
    assign process_intf_3.ap_start = AESL_inst_merge_sort.read_input_3_U0.ap_start;
    assign process_intf_3.ap_ready = AESL_inst_merge_sort.read_input_3_U0.ap_ready;
    assign process_intf_3.ap_done = AESL_inst_merge_sort.read_input_3_U0.ap_done;
    assign process_intf_3.ap_continue = AESL_inst_merge_sort.read_input_3_U0.ap_continue;
    assign process_intf_3.real_start = AESL_inst_merge_sort.read_input_3_U0.real_start;
    assign process_intf_3.pin_stall = 1'b0;
    assign process_intf_3.pout_stall = 1'b0 | ~AESL_inst_merge_sort.read_input_3_U0.right_stream_blk_n;
    assign process_intf_3.cin_stall = 1'b0;
    assign process_intf_3.cout_stall = 1'b0;
    assign process_intf_3.region_idle = region_0_idle;
    assign process_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_3;
    csv_file_dump pstatus_csv_dumper_3;
    df_process_monitor process_monitor_3;
    df_process_intf process_intf_4(clock,reset);
    assign process_intf_4.ap_start = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_start;
    assign process_intf_4.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_ready;
    assign process_intf_4.ap_done = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_done;
    assign process_intf_4.ap_continue = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_continue;
    assign process_intf_4.real_start = AESL_inst_merge_sort.merge_sort_iterative_1_U0.real_start;
    assign process_intf_4.pin_stall = 1'b0 | ~AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.left_stream_blk_n;
    assign process_intf_4.pout_stall = 1'b0 | ~AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.tmp_left_blk_n;
    assign process_intf_4.cin_stall = 1'b0;
    assign process_intf_4.cout_stall = 1'b0;
    assign process_intf_4.region_idle = region_0_idle;
    assign process_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_4;
    csv_file_dump pstatus_csv_dumper_4;
    df_process_monitor process_monitor_4;
    df_process_intf process_intf_5(clock,reset);
    assign process_intf_5.ap_start = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_start;
    assign process_intf_5.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_ready;
    assign process_intf_5.ap_done = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_done;
    assign process_intf_5.ap_continue = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_continue;
    assign process_intf_5.real_start = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_start;
    assign process_intf_5.pin_stall = 1'b0 | ~AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.right_stream_blk_n;
    assign process_intf_5.pout_stall = 1'b0 | ~AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.tmp_right_blk_n;
    assign process_intf_5.cin_stall = 1'b0;
    assign process_intf_5.cout_stall = 1'b0;
    assign process_intf_5.region_idle = region_0_idle;
    assign process_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_5;
    csv_file_dump pstatus_csv_dumper_5;
    df_process_monitor process_monitor_5;
    df_process_intf process_intf_6(clock,reset);
    assign process_intf_6.ap_start = AESL_inst_merge_sort.write_tmp_U0.ap_start;
    assign process_intf_6.ap_ready = AESL_inst_merge_sort.write_tmp_U0.ap_ready;
    assign process_intf_6.ap_done = AESL_inst_merge_sort.write_tmp_U0.ap_done;
    assign process_intf_6.ap_continue = AESL_inst_merge_sort.write_tmp_U0.ap_continue;
    assign process_intf_6.real_start = AESL_inst_merge_sort.write_tmp_U0.real_start;
    assign process_intf_6.pin_stall = 1'b0 | ~AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.tmp_right_blk_n | ~AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.tmp_left_blk_n;
    assign process_intf_6.pout_stall = 1'b0 | ~AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.tmp_blk_n | ~AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.tmp_blk_n;
    assign process_intf_6.cin_stall = 1'b0;
    assign process_intf_6.cout_stall = 1'b0;
    assign process_intf_6.region_idle = region_0_idle;
    assign process_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_6;
    csv_file_dump pstatus_csv_dumper_6;
    df_process_monitor process_monitor_6;
    df_process_intf process_intf_7(clock,reset);
    assign process_intf_7.ap_start = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_start;
    assign process_intf_7.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_ready;
    assign process_intf_7.ap_done = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_done;
    assign process_intf_7.ap_continue = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_continue;
    assign process_intf_7.real_start = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_start;
    assign process_intf_7.pin_stall = 1'b0 | ~AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.tmp_blk_n;
    assign process_intf_7.pout_stall = 1'b0 | ~AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.output_stream_blk_n;
    assign process_intf_7.cin_stall = 1'b0;
    assign process_intf_7.cout_stall = 1'b0;
    assign process_intf_7.region_idle = region_0_idle;
    assign process_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_7;
    csv_file_dump pstatus_csv_dumper_7;
    df_process_monitor process_monitor_7;
    df_process_intf process_intf_8(clock,reset);
    assign process_intf_8.ap_start = AESL_inst_merge_sort.write_output_U0.ap_start;
    assign process_intf_8.ap_ready = AESL_inst_merge_sort.write_output_U0.ap_ready;
    assign process_intf_8.ap_done = AESL_inst_merge_sort.write_output_U0.ap_done;
    assign process_intf_8.ap_continue = AESL_inst_merge_sort.write_output_U0.ap_continue;
    assign process_intf_8.real_start = AESL_inst_merge_sort.write_output_U0.ap_start;
    assign process_intf_8.pin_stall = 1'b0 | ~AESL_inst_merge_sort.write_output_U0.output_r_blk_n | ~AESL_inst_merge_sort.write_output_U0.output_stream_blk_n;
    assign process_intf_8.pout_stall = 1'b0;
    assign process_intf_8.cin_stall = 1'b0;
    assign process_intf_8.cout_stall = 1'b0;
    assign process_intf_8.region_idle = region_0_idle;
    assign process_intf_8.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_8;
    csv_file_dump pstatus_csv_dumper_8;
    df_process_monitor process_monitor_8;

    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_merge_sort.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_merge_sort.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_merge_sort.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_left_right_fu_4718.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_left_right_fu_4718.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_left_right_fu_4718.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_left_right_fu_4718.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_left_right_fu_4718.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_left_right_fu_4718.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_left_right_fu_5228.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_left_right_fu_5228.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_left_right_fu_5228.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;

    seq_loop_intf#(15) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_1.post_states_valid = 1'b1;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_ST_fsm_state13;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(15) seq_loop_monitor_1;
    seq_loop_intf#(15) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_2.pre_states_valid = 1'b1;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_ST_fsm_state14;
    assign seq_loop_intf_2.post_states_valid = 1'b1;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_2.quit_states_valid = 1'b1;
    assign seq_loop_intf_2.cur_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_merge_sort.merge_sort_iterative_1_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(15) seq_loop_monitor_2;
    seq_loop_intf#(15) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_3.pre_states_valid = 1'b1;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_3.post_states_valid = 1'b1;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_3.quit_states_valid = 1'b1;
    assign seq_loop_intf_3.cur_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_ST_fsm_state13;
    assign seq_loop_intf_3.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(15) seq_loop_monitor_3;
    seq_loop_intf#(15) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_4.pre_states_valid = 1'b1;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_ST_fsm_state14;
    assign seq_loop_intf_4.post_states_valid = 1'b1;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_4.quit_states_valid = 1'b1;
    assign seq_loop_intf_4.cur_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_merge_sort.merge_sort_iterative_2_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_4.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(15) seq_loop_monitor_4;
    seq_loop_intf#(15) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_5.pre_states_valid = 1'b1;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_5.post_states_valid = 1'b1;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_5.quit_states_valid = 1'b1;
    assign seq_loop_intf_5.cur_state = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_ST_fsm_state13;
    assign seq_loop_intf_5.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(15) seq_loop_monitor_5;
    seq_loop_intf#(15) seq_loop_intf_6(clock,reset);
    assign seq_loop_intf_6.pre_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_6.pre_states_valid = 1'b1;
    assign seq_loop_intf_6.post_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_ST_fsm_state14;
    assign seq_loop_intf_6.post_states_valid = 1'b1;
    assign seq_loop_intf_6.quit_loop_state0 = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_6.quit_states_valid = 1'b1;
    assign seq_loop_intf_6.cur_state = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_CS_fsm;
    assign seq_loop_intf_6.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_6.iter_end_state0 = AESL_inst_merge_sort.merge_sort_iterative_U0.ap_ST_fsm_state5;
    assign seq_loop_intf_6.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_6.one_state_loop = 1'b0;
    assign seq_loop_intf_6.one_state_block = 1'b0;
    assign seq_loop_intf_6.finish = finish;
    csv_file_dump seq_loop_csv_dumper_6;
    seq_loop_monitor #(15) seq_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_merge_sort.read_input_U0.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_merge_sort.read_input_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_merge_sort.read_input_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_merge_sort.read_input_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_merge_sort.read_input_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_merge_sort.read_input_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_merge_sort.read_input_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_merge_sort.read_input_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_merge_sort.read_input_U0.ap_enable_reg_pp0_iter10;
    assign upc_loop_intf_1.quit_enable = AESL_inst_merge_sort.read_input_U0.ap_enable_reg_pp0_iter10;
    assign upc_loop_intf_1.loop_start = AESL_inst_merge_sort.read_input_U0.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_merge_sort.read_input_U0.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_merge_sort.read_input_U0.ap_done;
    assign upc_loop_intf_1.loop_continue = AESL_inst_merge_sort.read_input_U0.ap_continue;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_merge_sort.read_input_3_U0.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_merge_sort.read_input_3_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_merge_sort.read_input_3_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_merge_sort.read_input_3_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_merge_sort.read_input_3_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_merge_sort.read_input_3_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_merge_sort.read_input_3_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_merge_sort.read_input_3_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_merge_sort.read_input_3_U0.ap_enable_reg_pp0_iter10;
    assign upc_loop_intf_2.quit_enable = AESL_inst_merge_sort.read_input_3_U0.ap_enable_reg_pp0_iter10;
    assign upc_loop_intf_2.loop_start = AESL_inst_merge_sort.read_input_3_U0.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_merge_sort.read_input_3_U0.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_merge_sort.read_input_3_U0.ap_done;
    assign upc_loop_intf_2.loop_continue = AESL_inst_merge_sort.read_input_3_U0.ap_continue;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(1) upc_loop_monitor_2;
    upc_loop_intf#(1) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.quit_enable = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.loop_start = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_fu_4200.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(1) upc_loop_monitor_3;
    upc_loop_intf#(1) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.quit_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_4.quit_enable = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_4.loop_start = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_merge_fu_5752.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(1) upc_loop_monitor_4;
    upc_loop_intf#(1) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.quit_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_5.quit_enable = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_5.loop_start = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_buffer_write_fu_5759.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b1;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(1) upc_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.quit_state = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.quit_enable = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.loop_start = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_merge_sort.merge_sort_iterative_1_U0.grp_merge_sort_iterative_1_Pipeline_output_fu_6791.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b1;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(1) upc_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.quit_enable = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.loop_start = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_fu_4200.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b1;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(1) upc_loop_monitor_7;
    upc_loop_intf#(1) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.quit_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_8.quit_enable = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_8.loop_start = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_merge_fu_5752.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b1;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(1) upc_loop_monitor_8;
    upc_loop_intf#(1) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_9.quit_enable = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_9.loop_start = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_buffer_write_fu_5759.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b1;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(1) upc_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.quit_enable = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.loop_start = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_merge_sort.merge_sort_iterative_2_U0.grp_merge_sort_iterative_2_Pipeline_output_fu_6791.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b1;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(1) upc_loop_monitor_10;
    upc_loop_intf#(1) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.quit_state = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.quit_enable = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.loop_start = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_108_1_fu_22.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b1;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(1) upc_loop_monitor_11;
    upc_loop_intf#(1) upc_loop_intf_12(clock,reset);
    assign upc_loop_intf_12.cur_state = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_CS_fsm;
    assign upc_loop_intf_12.iter_start_state = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_end_state = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.quit_state = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_start_block = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_end_block = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.quit_block = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_start_enable = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_12.iter_end_enable = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.quit_enable = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.loop_start = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_start;
    assign upc_loop_intf_12.loop_ready = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_ready;
    assign upc_loop_intf_12.loop_done = AESL_inst_merge_sort.write_tmp_U0.grp_write_tmp_Pipeline_VITIS_LOOP_113_2_fu_30.ap_done_int;
    assign upc_loop_intf_12.loop_continue = 1'b1;
    assign upc_loop_intf_12.quit_at_end = 1'b1;
    assign upc_loop_intf_12.finish = finish;
    csv_file_dump upc_loop_csv_dumper_12;
    upc_loop_monitor #(1) upc_loop_monitor_12;
    upc_loop_intf#(1) upc_loop_intf_13(clock,reset);
    assign upc_loop_intf_13.cur_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_CS_fsm;
    assign upc_loop_intf_13.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_end_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.quit_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_start_block = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_end_block = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.quit_block = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_start_enable = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_13.iter_end_enable = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.quit_enable = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.loop_start = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_start;
    assign upc_loop_intf_13.loop_ready = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_ready;
    assign upc_loop_intf_13.loop_done = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_fu_4198.ap_done_int;
    assign upc_loop_intf_13.loop_continue = 1'b1;
    assign upc_loop_intf_13.quit_at_end = 1'b1;
    assign upc_loop_intf_13.finish = finish;
    csv_file_dump upc_loop_csv_dumper_13;
    upc_loop_monitor #(1) upc_loop_monitor_13;
    upc_loop_intf#(1) upc_loop_intf_14(clock,reset);
    assign upc_loop_intf_14.cur_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_CS_fsm;
    assign upc_loop_intf_14.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_end_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.quit_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_start_block = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_end_block = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.quit_block = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_start_enable = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_14.iter_end_enable = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_14.quit_enable = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_14.loop_start = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_start;
    assign upc_loop_intf_14.loop_ready = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_ready;
    assign upc_loop_intf_14.loop_done = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_merge_fu_6262.ap_done_int;
    assign upc_loop_intf_14.loop_continue = 1'b1;
    assign upc_loop_intf_14.quit_at_end = 1'b1;
    assign upc_loop_intf_14.finish = finish;
    csv_file_dump upc_loop_csv_dumper_14;
    upc_loop_monitor #(1) upc_loop_monitor_14;
    upc_loop_intf#(1) upc_loop_intf_15(clock,reset);
    assign upc_loop_intf_15.cur_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_CS_fsm;
    assign upc_loop_intf_15.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_end_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.quit_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_start_block = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_end_block = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.quit_block = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_start_enable = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_15.iter_end_enable = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_15.quit_enable = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_15.loop_start = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_start;
    assign upc_loop_intf_15.loop_ready = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_ready;
    assign upc_loop_intf_15.loop_done = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_buffer_write_fu_6269.ap_done_int;
    assign upc_loop_intf_15.loop_continue = 1'b1;
    assign upc_loop_intf_15.quit_at_end = 1'b1;
    assign upc_loop_intf_15.finish = finish;
    csv_file_dump upc_loop_csv_dumper_15;
    upc_loop_monitor #(1) upc_loop_monitor_15;
    upc_loop_intf#(1) upc_loop_intf_16(clock,reset);
    assign upc_loop_intf_16.cur_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_CS_fsm;
    assign upc_loop_intf_16.iter_start_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_end_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.quit_state = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_start_block = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_end_block = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.quit_block = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_start_enable = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_16.iter_end_enable = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_16.quit_enable = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_16.loop_start = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_start;
    assign upc_loop_intf_16.loop_ready = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_ready;
    assign upc_loop_intf_16.loop_done = AESL_inst_merge_sort.merge_sort_iterative_U0.grp_merge_sort_iterative_Pipeline_output_fu_7301.ap_done_int;
    assign upc_loop_intf_16.loop_continue = 1'b1;
    assign upc_loop_intf_16.quit_at_end = 1'b1;
    assign upc_loop_intf_16.finish = finish;
    csv_file_dump upc_loop_csv_dumper_16;
    upc_loop_monitor #(1) upc_loop_monitor_16;
    upc_loop_intf#(1) upc_loop_intf_17(clock,reset);
    assign upc_loop_intf_17.cur_state = AESL_inst_merge_sort.write_output_U0.ap_CS_fsm;
    assign upc_loop_intf_17.iter_start_state = AESL_inst_merge_sort.write_output_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_end_state = AESL_inst_merge_sort.write_output_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.quit_state = AESL_inst_merge_sort.write_output_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_start_block = AESL_inst_merge_sort.write_output_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_end_block = AESL_inst_merge_sort.write_output_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.quit_block = AESL_inst_merge_sort.write_output_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_start_enable = AESL_inst_merge_sort.write_output_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_17.iter_end_enable = AESL_inst_merge_sort.write_output_U0.ap_enable_reg_pp0_iter8;
    assign upc_loop_intf_17.quit_enable = AESL_inst_merge_sort.write_output_U0.ap_enable_reg_pp0_iter8;
    assign upc_loop_intf_17.loop_start = AESL_inst_merge_sort.write_output_U0.ap_start;
    assign upc_loop_intf_17.loop_ready = AESL_inst_merge_sort.write_output_U0.ap_ready;
    assign upc_loop_intf_17.loop_done = AESL_inst_merge_sort.write_output_U0.ap_done;
    assign upc_loop_intf_17.loop_continue = AESL_inst_merge_sort.write_output_U0.ap_continue;
    assign upc_loop_intf_17.quit_at_end = 1'b1;
    assign upc_loop_intf_17.finish = finish;
    csv_file_dump upc_loop_csv_dumper_17;
    upc_loop_monitor #(1) upc_loop_monitor_17;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;

    fifo_csv_dumper_1 = new("./depth1.csv");
    cstatus_csv_dumper_1 = new("./chan_status1.csv");
    fifo_monitor_1 = new(fifo_csv_dumper_1,fifo_intf_1,cstatus_csv_dumper_1);
    fifo_csv_dumper_2 = new("./depth2.csv");
    cstatus_csv_dumper_2 = new("./chan_status2.csv");
    fifo_monitor_2 = new(fifo_csv_dumper_2,fifo_intf_2,cstatus_csv_dumper_2);
    fifo_csv_dumper_3 = new("./depth3.csv");
    cstatus_csv_dumper_3 = new("./chan_status3.csv");
    fifo_monitor_3 = new(fifo_csv_dumper_3,fifo_intf_3,cstatus_csv_dumper_3);
    fifo_csv_dumper_4 = new("./depth4.csv");
    cstatus_csv_dumper_4 = new("./chan_status4.csv");
    fifo_monitor_4 = new(fifo_csv_dumper_4,fifo_intf_4,cstatus_csv_dumper_4);
    fifo_csv_dumper_5 = new("./depth5.csv");
    cstatus_csv_dumper_5 = new("./chan_status5.csv");
    fifo_monitor_5 = new(fifo_csv_dumper_5,fifo_intf_5,cstatus_csv_dumper_5);
    fifo_csv_dumper_6 = new("./depth6.csv");
    cstatus_csv_dumper_6 = new("./chan_status6.csv");
    fifo_monitor_6 = new(fifo_csv_dumper_6,fifo_intf_6,cstatus_csv_dumper_6);
    fifo_csv_dumper_7 = new("./depth7.csv");
    cstatus_csv_dumper_7 = new("./chan_status7.csv");
    fifo_monitor_7 = new(fifo_csv_dumper_7,fifo_intf_7,cstatus_csv_dumper_7);

    pstall_csv_dumper_1 = new("./stalling1.csv");
    pstatus_csv_dumper_1 = new("./status1.csv");
    process_monitor_1 = new(pstall_csv_dumper_1,process_intf_1,pstatus_csv_dumper_1);
    pstall_csv_dumper_2 = new("./stalling2.csv");
    pstatus_csv_dumper_2 = new("./status2.csv");
    process_monitor_2 = new(pstall_csv_dumper_2,process_intf_2,pstatus_csv_dumper_2);
    pstall_csv_dumper_3 = new("./stalling3.csv");
    pstatus_csv_dumper_3 = new("./status3.csv");
    process_monitor_3 = new(pstall_csv_dumper_3,process_intf_3,pstatus_csv_dumper_3);
    pstall_csv_dumper_4 = new("./stalling4.csv");
    pstatus_csv_dumper_4 = new("./status4.csv");
    process_monitor_4 = new(pstall_csv_dumper_4,process_intf_4,pstatus_csv_dumper_4);
    pstall_csv_dumper_5 = new("./stalling5.csv");
    pstatus_csv_dumper_5 = new("./status5.csv");
    process_monitor_5 = new(pstall_csv_dumper_5,process_intf_5,pstatus_csv_dumper_5);
    pstall_csv_dumper_6 = new("./stalling6.csv");
    pstatus_csv_dumper_6 = new("./status6.csv");
    process_monitor_6 = new(pstall_csv_dumper_6,process_intf_6,pstatus_csv_dumper_6);
    pstall_csv_dumper_7 = new("./stalling7.csv");
    pstatus_csv_dumper_7 = new("./status7.csv");
    process_monitor_7 = new(pstall_csv_dumper_7,process_intf_7,pstatus_csv_dumper_7);
    pstall_csv_dumper_8 = new("./stalling8.csv");
    pstatus_csv_dumper_8 = new("./status8.csv");
    process_monitor_8 = new(pstall_csv_dumper_8,process_intf_8,pstatus_csv_dumper_8);

    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);



    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);
    seq_loop_csv_dumper_6 = new("./seq_loop_status6.csv");
    seq_loop_monitor_6 = new(seq_loop_intf_6,seq_loop_csv_dumper_6);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);
    upc_loop_csv_dumper_12 = new("./upc_loop_status12.csv");
    upc_loop_monitor_12 = new(upc_loop_intf_12,upc_loop_csv_dumper_12);
    upc_loop_csv_dumper_13 = new("./upc_loop_status13.csv");
    upc_loop_monitor_13 = new(upc_loop_intf_13,upc_loop_csv_dumper_13);
    upc_loop_csv_dumper_14 = new("./upc_loop_status14.csv");
    upc_loop_monitor_14 = new(upc_loop_intf_14,upc_loop_csv_dumper_14);
    upc_loop_csv_dumper_15 = new("./upc_loop_status15.csv");
    upc_loop_monitor_15 = new(upc_loop_intf_15,upc_loop_csv_dumper_15);
    upc_loop_csv_dumper_16 = new("./upc_loop_status16.csv");
    upc_loop_monitor_16 = new(upc_loop_intf_16,upc_loop_csv_dumper_16);
    upc_loop_csv_dumper_17 = new("./upc_loop_status17.csv");
    upc_loop_monitor_17 = new(upc_loop_intf_17,upc_loop_csv_dumper_17);

    sample_manager_inst.add_one_monitor(fifo_monitor_1);
    sample_manager_inst.add_one_monitor(fifo_monitor_2);
    sample_manager_inst.add_one_monitor(fifo_monitor_3);
    sample_manager_inst.add_one_monitor(fifo_monitor_4);
    sample_manager_inst.add_one_monitor(fifo_monitor_5);
    sample_manager_inst.add_one_monitor(fifo_monitor_6);
    sample_manager_inst.add_one_monitor(fifo_monitor_7);
    sample_manager_inst.add_one_monitor(process_monitor_1);
    sample_manager_inst.add_one_monitor(process_monitor_2);
    sample_manager_inst.add_one_monitor(process_monitor_3);
    sample_manager_inst.add_one_monitor(process_monitor_4);
    sample_manager_inst.add_one_monitor(process_monitor_5);
    sample_manager_inst.add_one_monitor(process_monitor_6);
    sample_manager_inst.add_one_monitor(process_monitor_7);
    sample_manager_inst.add_one_monitor(process_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_12);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_13);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_14);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_15);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_16);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_17);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1 || deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
